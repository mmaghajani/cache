library IEEE;
use IEEE.std_logic_1164.all;

entity lru_array is port (
  w1_select: out std_logic
  );
end lru_array;

architecture dataflow of lru_array is
begin

end dataflow;



