library IEEE;
use IEEE.std_logic_1164.all;

entity controller is port(
  write_request : in std_logic ;
  read_request: in std_logic ;
  ram_ready: in std_logic
  ) ;
end controller;

architecture behavioral of controller is
  constant s0: integer := 0 ;
  constant s0: integer := 0 ;
  constant s0: integer := 0 ;
  constant s0: integer := 0 ;
  
begin
  
end behavioral ;
